module ADDER_32B (
    input [31:0] in1,in2,
    output [31:0] out
    );

    assign out = in2 + in1;

endmodule