// tested and working perfect

module SIGN_EXTEND (
    input [15:0] in,
    output [31:0] out
);

assign out = in;

endmodule 